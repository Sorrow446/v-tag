module vtag