module tag