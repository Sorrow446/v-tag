module mp4

pub const (
	resolve_genre = {
		0x23: 'Acid'
		0x4B: 'Acid Jazz'
		0x4A: 'Acid Punk'
		0x64: 'Acoustic'
		0x15: 'Alternative'
		0x1B: 'Ambient'
		0x5B: 'Avantgarde'
		0x75: 'Ballad'
		0x2A: 'Bass'
		0x56: 'Bebob'
		0x61: 'Big Band'
		0x5A: 'Bluegrass'
		0x01: 'Blues'
		0x6C: 'Booty Bass'
		0x42: 'Cabaret'
		0x59: 'Celtic'
		0x69: 'Chamber Music'
		0x67: 'Chanson'
		0x62: 'Chorus'
		0x3E: 'Christian Rap'
		0x02: 'Classic Rock'
		0x21: 'Classical'
		0x71: 'Club'
		0x3A: 'Comedy'
		0x03: 'Country'
		0x3B: 'Cult'
		0x04: 'Dance'
		0x7E: 'Dance Hall'
		0x33: 'Darkwave'
		0x17: 'Death Metal'
		0x05: 'Disco'
		0x38: 'Dream'
		0x7B: 'Drum Solo'
		0x79: 'Duet'
		0x63: 'Easy Listening'
		0x35: 'Electronic'
		0x31: 'Ethnic'
		0x37: 'Eurodance'
		0x7D: 'Euro-House'
		0x1A: 'Euro-Techno'
		0x51: 'Folk'
		0x74: 'Folklore'
		0x78: 'Freestyle'
		0x06: 'Funk'
		0x1F: 'Fusion'
		0x25: 'Game'
		0x3C: 'Gangsta'
		0x27: 'Gospel'
		0x32: 'Gothic'
		0x5C: 'Gothic Rock'
		0x07: 'Grunge'
		0x50: 'Hard Rock'
		0x08: 'Hip-Hop'
		0x24: 'House'
		0x65: 'Humour'
		0x14: 'Industrial'
		0x22: 'Instrumental'
		0x2F: 'Instrumental Pop'
		0x30: 'Instrumental Rock'
		0x09: 'Jazz'
		0x1E: 'Jazz+Funk'
		0x40: 'Jungle'
		0x57: 'Latin'
		0x48: 'Lo-Fi'
		0x2E: 'Meditative'
		0x0A: 'Metal'
		0x4E: 'Musical'
		0x52: 'National Folk'
		0x41: 'Native American'
		0x0B: 'New Age'
		0x43: 'New Wave'
		0x28: 'Noise'
		0x0C: 'Oldies'
		0x68: 'Opera'
		0x0D: 'Other'
		0x4C: 'Polka'
		0x0E: 'Pop'
		0x3F: 'Pop/Funk'
		0x36: 'Pop-Folk'
		0x6E: 'Porn Groove'
		0x76: 'Power Ballad'
		0x18: 'Pranks'
		0x6D: 'Primus'
		0x5D: 'Progressive Rock'
		0x5E: 'Psychedelic Rock'
		0x2C: 'Punk'
		0x7A: 'Punk Rock'
		0x0F: 'R&B'
		0x10: 'Rap'
		0x45: 'Rave'
		0x11: 'Reggae'
		0x4D: 'Retro'
		0x58: 'Revival'
		0x77: 'Rhythmic Soul'
		0x12: 'Rock'
		0x4F: 'Rock & Roll'
		0x73: 'Samba'
		0x6F: 'Satire'
		0x46: 'Showtunes'
		0x16: 'Ska'
		0x70: 'Slow Jam'
		0x60: 'Slow Rock'
		0x6A: 'Sonata'
		0x2B: 'Soul'
		0x26: 'Sound Clip'
		0x19: 'Soundtrack'
		0x39: 'Southern Rock'
		0x2D: 'Space'
		0x66: 'Speech'
		0x54: 'Swing'
		0x5F: 'Symphonic Rock'
		0x6B: 'Symphony'
		0x72: 'Tango'
		0x13: 'Techno'
		0x34: 'Techno-Industrial'
		0x3D: 'Top 40'
		0x47: 'Trailer'
		0x20: 'Trance'
		0x49: 'Tribal'
		0x1C: 'Trip-Hop'
		0x1D: 'Vocal'
	}

	resolve_atom = {
		'a9616c62': 'album'
		'61415254': 'album_artist'
		'736f6161': 'album_artist_sort'
		'736f616c': 'album_sort'
		'a9415254': 'artist'
		'736f6172': 'artist_sort'
		//'746d706f': 'bpm',
		'a9636d74': 'comment'
		'a9777274': 'composer'
		'736f636f': 'composer_sort'
		//'6370696c': 'compilation',
		'a9636f6e': 'conductor'
		'63707274': 'copyright'
		'a967656e': 'genre'
		//'676e7265': 'genre',
		'6f776e72': 'owner'
		'74766573': 'tv_episode'
		'64657363': 'description'
		'a9746f6f': 'encoder'
		'a96e7274': 'narrator'
		//'70637374': 'podcast',
		'a9707562': 'publisher'
		// '63617467': 'podcast_category',
		// '6c646573': 'podcast_description',
		// '6b657977': 'podcast_keywords',
		// '7075726c': 'podcast_url',
		'a96e616d': 'title'
		'736f6e6d': 'title_sort'
		'736f736e': 'tv_show_sort'
		'a96c7972': 'unsynced_lyrics'
		'a9646179': 'year'
		// egid, int
		//'65676964': 'podcast_id',
		// ©mvc, int
		//'a96d7663': 'movement_total'
	}

	nums = [48, 49, 50, 51, 52, 53, 54, 55, 56, 57]
)
