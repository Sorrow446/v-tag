module tag

pub const (
	resolve_field_flac = {
		'album': 'album',
		'albumartist': 'album_artist',
		'artist': 'artist',
		'comment': 'comment',
		'contact': 'contact',
		'copyright': 'copyright',
		'date': 'date',
		'encoder': 'encoder',
		'genre': 'genre',
		'isrc': 'isrc',
		'itunesadvisory': 'itunes_advisory',
		'label': 'label',
		'performer': 'performer',
		'publisher': 'publisher',
		'title': 'title',
	}

	resolve_field_id3 = {
		'TPE2': 'album_artist'
		'TALB': 'album',
		'TPE1': 'artist',
		'TCON': 'genre',
		'COMM': 'comment',
		'TIT2': 'title',
		'TCOP': 'copyright',
		'TCOM': 'composer',
		'TPE3': 'conductor',
		'TENC': 'encoded_by',
		'TIT1': 'content_group',
		'TSRC': 'isrc',
		'TPUB': 'publisher',
		'WXXX': 'www',
		'USLT': 'unsynced_lyrics',
		'TDAT': 'date',
	}

	resolve_pic_type_flac = {
		0: 'Other',
		1: 'Icon',
		2: 'Other Icon',
		3: 'Front Cover',
		4: 'Back Cover',
		5: 'Leaflet',
		6: 'Media',
		7: 'Lead Artist',
		8: 'Artist',
		9: 'Conductor',
		10: 'Band',
		11: 'Composer',
		12: 'Lyricist',
		13: 'Recording Location',
		14: 'During Recording',
		15: 'During Performance',
		16: 'Video Capture',
		18: 'Illustration',
		19: 'Band Logotype',
		20: 'Publisher Logotype',
	}

	resolve_pic_type_id3 = {
		0x0:  'Other',
		0x01: 'Icon',
		0x02: 'Other Icon',
		0x03: 'Front Cover',
		0x04: 'Back Cover',
		0x05: 'Leaflet',
		0x06: 'Media',
		0x07: 'Lead Artist',
		0x08: 'Artist',
		0x09: 'Conductor',
		0x0A: 'Band',
		0x0B: 'Composer',
		0x0C: 'Lyricist',
		0x0D: 'Recording Location',
		0x0E: 'During Recording',
		0x0F: 'During Performance',
		0x1:  'Video Capture',
		0x12: 'Illustration',
		0x13: 'Band Logotype',
		0x14: 'Publisher Logotype',
	}

	id3_frames = [
		'TPE2', 'TALB', 'TPE1', 'TCON',
		'COMM', 'TIT2', 'TCOP', 'TCOM',
		'TENC', 'TXXX', 'TRCK', 'TPOS',
		'TYER', 'TBPM', 'TBMP', 'TCMP',
		'TPE3', 'TIT1', 'TSRC', 'TPUB',
		'WXXX', 'USLT', 'TDAT', 'APIC',
	]

	resolve_genre = {
		'(0)': 'Blues',
	  	'(1)': 'Classic Rock',
	  	'(2)': 'Country',
	  	'(3)': 'Dance',
	  	'(4)': 'Disco',
	  	'(5)': 'Funk',
	  	'(6)': 'Grunge',
	  	'(7)': 'Hip-Hop',
	  	'(8)': 'Jazz',
	  	'(9)': 'Metal',
	  	'(10)': 'New Age',
	  	'(11)': 'Oldies',
		'(12)': 'Other',
		'(13)': 'Pop',
		'(14)': 'R&B',
		'(15)': 'Rap',
		'(16)': 'Reggae',
		'(17)': 'Rock',
		'(18)': 'Techno',
		'(19)': 'Industrial',
		'(20)': 'Alternative',
		'(21)': 'Ska',
		'(22)': 'Death Metal',
		'(23)': 'Pranks',
		'(24)': 'Soundtrack',
		'(25)': 'Euro-Techno',
		'(26)': 'Ambient',
		'(27)': 'Trip-Hop',
		'(28)': 'Vocal',
		'(29)': 'Jazz+Funk',
		'(30)': 'Fusion',
		'(31)': 'Trance',
		'(32)': 'Classical',
		'(33)': 'Instrumental',
		'(34)': 'Acid',
		'(35)': 'House',
		'(36)': 'Game',
		'(37)': 'Sound Clip',
		'(38)': 'Gospel',
		'(39)': 'Noise',
		'(40)': 'AlternRock',
		'(41)': 'Bass',
		'(42)': 'Soul',
		'(43)': 'Punk',
		'(44)': 'Space',
		'(45)': 'Meditative',
		'(46)': 'Instrumental Pop',
		'(47)': 'Instrumental Rock',
		'(48)': 'Ethnic',
		'(49)': 'Gothic',
		'(50)': 'Darkwave',
		'(51)': 'Techno-Industrial',
		'(52)': 'Electronic',
		'(53)': 'Pop-Folk',
		'(54)': 'Eurodance',
		'(55)': 'Dream',
		'(56)': 'Southern Rock',
		'(57)': 'Comedy',
		'(58)': 'Cult',
		'(59)': 'Gangsta',
		'(60)': 'Top 40',
		'(61)': 'Christian Rap',
		'(62)': 'Pop/Funk',
		'(63)': 'Jungle',
		'(64)': 'Native American',
		'(65)': 'Cabaret',
		'(66)': 'New Wave',
		'(67)': 'Psychadelic',
		'(68)': 'Rave',
		'(69)': 'Showtunes',
		'(70)': 'Trailer',
		'(71)': 'Lo-Fi',
		'(72)': 'Tribal',
		'(73)': 'Acid Punk',
		'(74)': 'Acid Jazz',
		'(75)': 'Polka',
		'(76)': 'Retro',
		'(77)': 'Musical',
		'(78)': 'Rock & Roll',
		'(79)': 'Hard Rock',
		'(80)': 'Folk',
		'(81)': 'Folk-Rock',
		'(82)': 'National Folk',
		'(83)': 'Swing',
		'(84)': 'Fast Fusion',
		'(85)': 'Bebob',
		'(86)': 'Latin',
		'(87)': 'Revival',
		'(88)': 'Celtic',
		'(89)': 'Bluegrass',
		'(90)': 'Avantgarde',
		'(91)': 'Gothic Rock',
		'(92)': 'Progressive Rock',
		'(93)': 'Psychedelic Rock',
		'(94)': 'Symphonic Rock',
		'(95)': 'Slow Rock',
		'(96)': 'Big Band',
		'(97)': 'Chorus',
		'(98)': 'Easy Listening',
		'(99)': 'Acoustic',
		'(100)': 'Humour',
		'(101)': 'Speech',
		'(102)': 'Chanson',
		'(103)': 'Opera',
		'(104)': 'Chamber Music',
		'(105)': 'Sonata',
		'(106)': 'Symphony',
		'(107)': 'Booty Bass',
		'(108)': 'Primus',
		'(109)': 'Porn Groove',
		'(110)': 'Satire',
		'(111)': 'Slow Jam',
		'(112)': 'Club',
		'(113)': 'Tango',
		'(114)': 'Samba',
		'(115)': 'Folklore',
		'(116)': 'Ballad',
		'(117)': 'Power Ballad',
		'(118)': 'Rhythmic Soul',
		'(119)': 'Freestyle',
		'(120)': 'Duet',
		'(121)': 'Punk Rock',
		'(122)': 'Drum Solo',
		'(123)': 'A cappella',
		'(124)': 'Euro-House',
		'(125)': 'Dance Hall',
	}
)